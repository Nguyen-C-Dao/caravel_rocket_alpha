VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper1
  CLASS BLOCK ;
  FOREIGN user_project_wrapper1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2880.000 BY 3480.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1410.740 2884.800 1411.940 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2199.210 3479.000 2199.770 3484.800 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1879.510 3479.000 1880.070 3484.800 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1559.350 3479.000 1559.910 3484.800 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.190 3479.000 1239.750 3484.800 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.490 3479.000 920.050 3484.800 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.330 3479.000 599.890 3484.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.170 3479.000 279.730 3484.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3447.340 1.000 3448.540 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3189.620 1.000 3190.820 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2931.900 1.000 2933.100 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1673.900 2884.800 1675.100 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2673.500 1.000 2674.700 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2415.780 1.000 2416.980 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2158.060 1.000 2159.260 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1900.340 1.000 1901.540 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1642.620 1.000 1643.820 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1384.900 1.000 1386.100 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1127.180 1.000 1128.380 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 869.460 1.000 870.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 611.740 1.000 612.940 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1936.380 2884.800 1937.580 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2198.860 2884.800 2200.060 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2461.340 2884.800 2462.540 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2724.500 2884.800 2725.700 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2986.980 2884.800 2988.180 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 3249.460 2884.800 3250.660 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2839.530 3479.000 2840.090 3484.800 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2519.370 3479.000 2519.930 3484.800 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 32.380 2884.800 33.580 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2264.820 2884.800 2266.020 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2527.300 2884.800 2528.500 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2789.780 2884.800 2790.980 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 3052.940 2884.800 3054.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 3315.420 2884.800 3316.620 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2759.490 3479.000 2760.050 3484.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2439.330 3479.000 2439.890 3484.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2119.170 3479.000 2119.730 3484.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.470 3479.000 1800.030 3484.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1479.310 3479.000 1479.870 3484.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 228.900 2884.800 230.100 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.150 3479.000 1159.710 3484.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.450 3479.000 840.010 3484.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.290 3479.000 519.850 3484.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.130 3479.000 199.690 3484.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3382.740 1.000 3383.940 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3125.020 1.000 3126.220 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2867.300 1.000 2868.500 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2609.580 1.000 2610.780 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2351.860 1.000 2353.060 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2093.460 1.000 2094.660 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 426.100 2884.800 427.300 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1835.740 1.000 1836.940 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1578.020 1.000 1579.220 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1320.300 1.000 1321.500 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1062.580 1.000 1063.780 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 804.860 1.000 806.060 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 547.140 1.000 548.340 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 353.340 1.000 354.540 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 160.220 1.000 161.420 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 623.300 2884.800 624.500 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 819.820 2884.800 821.020 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1017.020 2884.800 1018.220 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1214.220 2884.800 1215.420 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1476.700 2884.800 1477.900 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1739.180 2884.800 1740.380 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2001.660 2884.800 2002.860 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 163.620 2884.800 164.820 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2396.060 2884.800 2397.260 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2658.540 2884.800 2659.740 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2921.020 2884.800 2922.220 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 3184.180 2884.800 3185.380 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 3446.660 2884.800 3447.860 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2599.410 3479.000 2599.970 3484.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2279.250 3479.000 2279.810 3484.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.550 3479.000 1960.110 3484.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.390 3479.000 1639.950 3484.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1319.230 3479.000 1319.790 3484.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 360.140 2884.800 361.340 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.530 3479.000 1000.090 3484.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.370 3479.000 679.930 3484.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.210 3479.000 359.770 3484.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.510 3479.000 40.070 3484.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3253.540 1.000 3254.740 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2995.820 1.000 2997.020 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2738.100 1.000 2739.300 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2480.380 1.000 2481.580 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2222.660 1.000 2223.860 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1964.940 1.000 1966.140 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 557.340 2884.800 558.540 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1707.220 1.000 1708.420 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1449.500 1.000 1450.700 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1191.780 1.000 1192.980 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 933.380 1.000 934.580 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 675.660 1.000 676.860 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 417.940 1.000 419.140 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 224.820 1.000 226.020 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 31.700 1.000 32.900 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 754.540 2884.800 755.740 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 951.060 2884.800 952.260 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1148.260 2884.800 1149.460 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1345.460 2884.800 1346.660 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1607.940 2884.800 1609.140 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1870.420 2884.800 1871.620 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2133.580 2884.800 2134.780 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 97.660 2884.800 98.860 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2330.100 2884.800 2331.300 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2593.260 2884.800 2594.460 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2855.740 2884.800 2856.940 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 3118.220 2884.800 3119.420 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 3380.700 2884.800 3381.900 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2679.450 3479.000 2680.010 3484.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2359.290 3479.000 2359.850 3484.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2039.130 3479.000 2039.690 3484.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1719.430 3479.000 1719.990 3484.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1399.270 3479.000 1399.830 3484.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 294.860 2884.800 296.060 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.110 3479.000 1079.670 3484.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.410 3479.000 759.970 3484.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.250 3479.000 439.810 3484.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.090 3479.000 119.650 3484.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3318.140 1.000 3319.340 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3060.420 1.000 3061.620 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2802.700 1.000 2803.900 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2544.980 1.000 2546.180 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2287.260 1.000 2288.460 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2029.540 1.000 2030.740 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 491.380 2884.800 492.580 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1771.820 1.000 1773.020 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1513.420 1.000 1514.620 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1255.700 1.000 1256.900 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 997.980 1.000 999.180 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 740.260 1.000 741.460 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 482.540 1.000 483.740 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 289.420 1.000 290.620 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 95.620 1.000 96.820 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 688.580 2884.800 689.780 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 885.780 2884.800 886.980 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1082.980 2884.800 1084.180 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1279.500 2884.800 1280.700 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1542.660 2884.800 1543.860 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1805.140 2884.800 1806.340 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2067.620 2884.800 2068.820 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.490 -4.800 621.050 1.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2369.410 -4.800 2369.970 1.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2386.890 -4.800 2387.450 1.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2404.370 -4.800 2404.930 1.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2421.850 -4.800 2422.410 1.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2439.330 -4.800 2439.890 1.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2456.810 -4.800 2457.370 1.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2474.290 -4.800 2474.850 1.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2491.770 -4.800 2492.330 1.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2509.250 -4.800 2509.810 1.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2526.730 -4.800 2527.290 1.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.290 -4.800 795.850 1.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2544.210 -4.800 2544.770 1.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2561.690 -4.800 2562.250 1.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2579.170 -4.800 2579.730 1.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2596.650 -4.800 2597.210 1.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2614.130 -4.800 2614.690 1.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2632.070 -4.800 2632.630 1.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2649.550 -4.800 2650.110 1.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2667.030 -4.800 2667.590 1.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2684.510 -4.800 2685.070 1.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2701.990 -4.800 2702.550 1.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.770 -4.800 813.330 1.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2719.470 -4.800 2720.030 1.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2736.950 -4.800 2737.510 1.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2754.430 -4.800 2754.990 1.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2771.910 -4.800 2772.470 1.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2789.390 -4.800 2789.950 1.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2806.870 -4.800 2807.430 1.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2824.350 -4.800 2824.910 1.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2841.830 -4.800 2842.390 1.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.250 -4.800 830.810 1.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.730 -4.800 848.290 1.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.210 -4.800 865.770 1.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.690 -4.800 883.250 1.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.170 -4.800 900.730 1.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.650 -4.800 918.210 1.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.130 -4.800 935.690 1.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.610 -4.800 953.170 1.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.970 -4.800 638.530 1.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.090 -4.800 970.650 1.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.570 -4.800 988.130 1.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.050 -4.800 1005.610 1.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.530 -4.800 1023.090 1.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.010 -4.800 1040.570 1.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1057.950 -4.800 1058.510 1.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.430 -4.800 1075.990 1.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.910 -4.800 1093.470 1.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.390 -4.800 1110.950 1.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.870 -4.800 1128.430 1.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.450 -4.800 656.010 1.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.350 -4.800 1145.910 1.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.830 -4.800 1163.390 1.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1180.310 -4.800 1180.870 1.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.790 -4.800 1198.350 1.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1215.270 -4.800 1215.830 1.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1232.750 -4.800 1233.310 1.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1250.230 -4.800 1250.790 1.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1267.710 -4.800 1268.270 1.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.190 -4.800 1285.750 1.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1302.670 -4.800 1303.230 1.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.930 -4.800 673.490 1.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.150 -4.800 1320.710 1.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1337.630 -4.800 1338.190 1.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.110 -4.800 1355.670 1.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1372.590 -4.800 1373.150 1.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1390.070 -4.800 1390.630 1.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.550 -4.800 1408.110 1.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1425.030 -4.800 1425.590 1.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1442.510 -4.800 1443.070 1.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1459.990 -4.800 1460.550 1.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1477.470 -4.800 1478.030 1.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.410 -4.800 690.970 1.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.950 -4.800 1495.510 1.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1512.430 -4.800 1512.990 1.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1529.910 -4.800 1530.470 1.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1547.390 -4.800 1547.950 1.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1564.870 -4.800 1565.430 1.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1582.350 -4.800 1582.910 1.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1599.830 -4.800 1600.390 1.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1617.310 -4.800 1617.870 1.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1634.790 -4.800 1635.350 1.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1652.270 -4.800 1652.830 1.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.890 -4.800 708.450 1.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1669.750 -4.800 1670.310 1.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.230 -4.800 1687.790 1.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.710 -4.800 1705.270 1.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.190 -4.800 1722.750 1.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1739.670 -4.800 1740.230 1.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1757.150 -4.800 1757.710 1.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1774.630 -4.800 1775.190 1.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1792.110 -4.800 1792.670 1.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1809.590 -4.800 1810.150 1.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1827.070 -4.800 1827.630 1.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.370 -4.800 725.930 1.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.010 -4.800 1845.570 1.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1862.490 -4.800 1863.050 1.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1879.970 -4.800 1880.530 1.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1897.450 -4.800 1898.010 1.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1914.930 -4.800 1915.490 1.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1932.410 -4.800 1932.970 1.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1949.890 -4.800 1950.450 1.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1967.370 -4.800 1967.930 1.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1984.850 -4.800 1985.410 1.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2002.330 -4.800 2002.890 1.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.850 -4.800 743.410 1.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2019.810 -4.800 2020.370 1.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2037.290 -4.800 2037.850 1.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2054.770 -4.800 2055.330 1.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2072.250 -4.800 2072.810 1.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.730 -4.800 2090.290 1.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2107.210 -4.800 2107.770 1.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2124.690 -4.800 2125.250 1.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2142.170 -4.800 2142.730 1.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2159.650 -4.800 2160.210 1.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2177.130 -4.800 2177.690 1.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.330 -4.800 760.890 1.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2194.610 -4.800 2195.170 1.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2212.090 -4.800 2212.650 1.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2229.570 -4.800 2230.130 1.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2247.050 -4.800 2247.610 1.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2264.530 -4.800 2265.090 1.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2282.010 -4.800 2282.570 1.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2299.490 -4.800 2300.050 1.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2316.970 -4.800 2317.530 1.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2334.450 -4.800 2335.010 1.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2351.930 -4.800 2352.490 1.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.810 -4.800 778.370 1.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.470 -4.800 627.030 1.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2375.390 -4.800 2375.950 1.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.870 -4.800 2393.430 1.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2410.350 -4.800 2410.910 1.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2427.830 -4.800 2428.390 1.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2445.310 -4.800 2445.870 1.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2462.790 -4.800 2463.350 1.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2480.270 -4.800 2480.830 1.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2497.750 -4.800 2498.310 1.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2515.230 -4.800 2515.790 1.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2532.710 -4.800 2533.270 1.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.270 -4.800 801.830 1.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2550.190 -4.800 2550.750 1.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2567.670 -4.800 2568.230 1.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2585.150 -4.800 2585.710 1.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2602.630 -4.800 2603.190 1.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2620.110 -4.800 2620.670 1.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2637.590 -4.800 2638.150 1.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2655.070 -4.800 2655.630 1.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2672.550 -4.800 2673.110 1.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2690.030 -4.800 2690.590 1.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2707.510 -4.800 2708.070 1.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.750 -4.800 819.310 1.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2724.990 -4.800 2725.550 1.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2742.470 -4.800 2743.030 1.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2759.950 -4.800 2760.510 1.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2777.430 -4.800 2777.990 1.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2794.910 -4.800 2795.470 1.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2812.390 -4.800 2812.950 1.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2829.870 -4.800 2830.430 1.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2847.350 -4.800 2847.910 1.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 836.230 -4.800 836.790 1.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.710 -4.800 854.270 1.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.190 -4.800 871.750 1.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.670 -4.800 889.230 1.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.150 -4.800 906.710 1.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.630 -4.800 924.190 1.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.110 -4.800 941.670 1.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.590 -4.800 959.150 1.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.950 -4.800 644.510 1.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.070 -4.800 976.630 1.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.550 -4.800 994.110 1.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.030 -4.800 1011.590 1.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1028.510 -4.800 1029.070 1.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1045.990 -4.800 1046.550 1.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1063.470 -4.800 1064.030 1.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.950 -4.800 1081.510 1.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.430 -4.800 1098.990 1.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1115.910 -4.800 1116.470 1.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.390 -4.800 1133.950 1.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.430 -4.800 661.990 1.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.870 -4.800 1151.430 1.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.350 -4.800 1168.910 1.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.830 -4.800 1186.390 1.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1203.310 -4.800 1203.870 1.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.790 -4.800 1221.350 1.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1238.270 -4.800 1238.830 1.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.750 -4.800 1256.310 1.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.230 -4.800 1273.790 1.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1290.710 -4.800 1291.270 1.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.190 -4.800 1308.750 1.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.910 -4.800 679.470 1.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.130 -4.800 1326.690 1.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1343.610 -4.800 1344.170 1.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1361.090 -4.800 1361.650 1.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.570 -4.800 1379.130 1.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1396.050 -4.800 1396.610 1.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.530 -4.800 1414.090 1.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1431.010 -4.800 1431.570 1.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1448.490 -4.800 1449.050 1.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.970 -4.800 1466.530 1.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1483.450 -4.800 1484.010 1.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.390 -4.800 696.950 1.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.930 -4.800 1501.490 1.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1518.410 -4.800 1518.970 1.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1535.890 -4.800 1536.450 1.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1553.370 -4.800 1553.930 1.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1570.850 -4.800 1571.410 1.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.330 -4.800 1588.890 1.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1605.810 -4.800 1606.370 1.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1623.290 -4.800 1623.850 1.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1640.770 -4.800 1641.330 1.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.250 -4.800 1658.810 1.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.870 -4.800 714.430 1.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.730 -4.800 1676.290 1.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.210 -4.800 1693.770 1.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.690 -4.800 1711.250 1.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.170 -4.800 1728.730 1.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1745.650 -4.800 1746.210 1.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1763.130 -4.800 1763.690 1.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1780.610 -4.800 1781.170 1.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1798.090 -4.800 1798.650 1.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1815.570 -4.800 1816.130 1.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1833.050 -4.800 1833.610 1.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.350 -4.800 731.910 1.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1850.530 -4.800 1851.090 1.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1868.010 -4.800 1868.570 1.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1885.490 -4.800 1886.050 1.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1902.970 -4.800 1903.530 1.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1920.450 -4.800 1921.010 1.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1937.930 -4.800 1938.490 1.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1955.410 -4.800 1955.970 1.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1972.890 -4.800 1973.450 1.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1990.370 -4.800 1990.930 1.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2007.850 -4.800 2008.410 1.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.830 -4.800 749.390 1.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2025.330 -4.800 2025.890 1.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2042.810 -4.800 2043.370 1.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2060.290 -4.800 2060.850 1.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2077.770 -4.800 2078.330 1.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2095.250 -4.800 2095.810 1.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2113.190 -4.800 2113.750 1.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.670 -4.800 2131.230 1.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2148.150 -4.800 2148.710 1.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2165.630 -4.800 2166.190 1.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.110 -4.800 2183.670 1.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.310 -4.800 766.870 1.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2200.590 -4.800 2201.150 1.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.070 -4.800 2218.630 1.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2235.550 -4.800 2236.110 1.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2253.030 -4.800 2253.590 1.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2270.510 -4.800 2271.070 1.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2287.990 -4.800 2288.550 1.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2305.470 -4.800 2306.030 1.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2322.950 -4.800 2323.510 1.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2340.430 -4.800 2340.990 1.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2357.910 -4.800 2358.470 1.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.790 -4.800 784.350 1.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.990 -4.800 632.550 1.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2381.370 -4.800 2381.930 1.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2398.850 -4.800 2399.410 1.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2416.330 -4.800 2416.890 1.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2433.810 -4.800 2434.370 1.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2451.290 -4.800 2451.850 1.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2468.770 -4.800 2469.330 1.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2486.250 -4.800 2486.810 1.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2503.730 -4.800 2504.290 1.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2521.210 -4.800 2521.770 1.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2538.690 -4.800 2539.250 1.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.250 -4.800 807.810 1.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2556.170 -4.800 2556.730 1.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2573.650 -4.800 2574.210 1.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2591.130 -4.800 2591.690 1.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2608.610 -4.800 2609.170 1.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2626.090 -4.800 2626.650 1.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2643.570 -4.800 2644.130 1.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2661.050 -4.800 2661.610 1.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2678.530 -4.800 2679.090 1.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2696.010 -4.800 2696.570 1.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2713.490 -4.800 2714.050 1.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.730 -4.800 825.290 1.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2730.970 -4.800 2731.530 1.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2748.450 -4.800 2749.010 1.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2765.930 -4.800 2766.490 1.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2783.410 -4.800 2783.970 1.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2800.890 -4.800 2801.450 1.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2818.370 -4.800 2818.930 1.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2835.850 -4.800 2836.410 1.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2853.330 -4.800 2853.890 1.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.210 -4.800 842.770 1.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.690 -4.800 860.250 1.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.170 -4.800 877.730 1.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.650 -4.800 895.210 1.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.130 -4.800 912.690 1.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.610 -4.800 930.170 1.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.090 -4.800 947.650 1.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 964.570 -4.800 965.130 1.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.470 -4.800 650.030 1.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.050 -4.800 982.610 1.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.530 -4.800 1000.090 1.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.010 -4.800 1017.570 1.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1034.490 -4.800 1035.050 1.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.970 -4.800 1052.530 1.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.450 -4.800 1070.010 1.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.930 -4.800 1087.490 1.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.410 -4.800 1104.970 1.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.890 -4.800 1122.450 1.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.370 -4.800 1139.930 1.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.950 -4.800 667.510 1.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.850 -4.800 1157.410 1.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.330 -4.800 1174.890 1.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.810 -4.800 1192.370 1.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1209.290 -4.800 1209.850 1.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.770 -4.800 1227.330 1.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1244.250 -4.800 1244.810 1.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.730 -4.800 1262.290 1.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.210 -4.800 1279.770 1.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1296.690 -4.800 1297.250 1.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.170 -4.800 1314.730 1.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.430 -4.800 684.990 1.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1331.650 -4.800 1332.210 1.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.130 -4.800 1349.690 1.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1366.610 -4.800 1367.170 1.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1384.090 -4.800 1384.650 1.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1401.570 -4.800 1402.130 1.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.050 -4.800 1419.610 1.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.530 -4.800 1437.090 1.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1454.010 -4.800 1454.570 1.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.490 -4.800 1472.050 1.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1488.970 -4.800 1489.530 1.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.910 -4.800 702.470 1.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1506.450 -4.800 1507.010 1.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.930 -4.800 1524.490 1.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1541.410 -4.800 1541.970 1.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1558.890 -4.800 1559.450 1.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1576.830 -4.800 1577.390 1.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1594.310 -4.800 1594.870 1.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1611.790 -4.800 1612.350 1.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1629.270 -4.800 1629.830 1.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1646.750 -4.800 1647.310 1.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1664.230 -4.800 1664.790 1.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.390 -4.800 719.950 1.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1681.710 -4.800 1682.270 1.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.190 -4.800 1699.750 1.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.670 -4.800 1717.230 1.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1734.150 -4.800 1734.710 1.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.630 -4.800 1752.190 1.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1769.110 -4.800 1769.670 1.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1786.590 -4.800 1787.150 1.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1804.070 -4.800 1804.630 1.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1821.550 -4.800 1822.110 1.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1839.030 -4.800 1839.590 1.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.870 -4.800 737.430 1.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1856.510 -4.800 1857.070 1.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1873.990 -4.800 1874.550 1.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1891.470 -4.800 1892.030 1.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1908.950 -4.800 1909.510 1.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1926.430 -4.800 1926.990 1.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1943.910 -4.800 1944.470 1.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1961.390 -4.800 1961.950 1.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1978.870 -4.800 1979.430 1.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1996.350 -4.800 1996.910 1.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2013.830 -4.800 2014.390 1.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.350 -4.800 754.910 1.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2031.310 -4.800 2031.870 1.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.790 -4.800 2049.350 1.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2066.270 -4.800 2066.830 1.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2083.750 -4.800 2084.310 1.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2101.230 -4.800 2101.790 1.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.710 -4.800 2119.270 1.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2136.190 -4.800 2136.750 1.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2153.670 -4.800 2154.230 1.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2171.150 -4.800 2171.710 1.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2188.630 -4.800 2189.190 1.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.830 -4.800 772.390 1.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2206.110 -4.800 2206.670 1.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2223.590 -4.800 2224.150 1.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2241.070 -4.800 2241.630 1.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2258.550 -4.800 2259.110 1.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2276.030 -4.800 2276.590 1.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2293.510 -4.800 2294.070 1.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2310.990 -4.800 2311.550 1.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2328.470 -4.800 2329.030 1.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2345.950 -4.800 2346.510 1.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2363.890 -4.800 2364.450 1.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.770 -4.800 790.330 1.000 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2859.310 -4.800 2859.870 1.000 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2864.830 -4.800 2865.390 1.000 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2870.810 -4.800 2871.370 1.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2876.790 -4.800 2877.350 1.000 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 14.090 2874.080 17.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 194.090 2874.080 197.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 374.090 2874.080 377.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 554.090 2874.080 557.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 734.090 2874.080 737.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 914.090 2874.080 917.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 1094.090 2874.080 1097.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 1274.090 2874.080 1277.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 1454.090 2874.080 1457.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 1634.090 2874.080 1637.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 1814.090 2874.080 1817.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 1994.090 2874.080 1997.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 2174.090 2874.080 2177.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 2354.090 2874.080 2357.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 2534.090 2874.080 2537.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 2714.090 2874.080 2717.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 2894.090 2874.080 2897.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 3074.090 2874.080 3077.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 3254.090 2874.080 3257.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 3434.090 2874.080 3437.190 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 10.640 192.070 240.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 10.640 372.070 240.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 10.640 552.070 240.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 10.640 732.070 240.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 10.640 2172.070 240.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 10.640 2352.070 240.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 10.640 2532.070 240.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 10.640 2712.070 240.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2802.470 241.840 2805.570 672.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 676.300 192.070 790.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 676.300 372.070 790.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 676.300 552.070 790.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 676.300 732.070 790.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 676.300 2172.070 790.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 676.300 2352.070 790.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 676.300 2532.070 790.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 676.300 2712.070 790.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2802.470 791.280 2805.570 1221.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 1226.300 192.070 1340.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 1226.300 372.070 1340.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 1226.300 552.070 1340.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 1226.300 732.070 1340.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 1226.300 2172.070 1340.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 1226.300 2352.070 1340.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 1226.300 2532.070 1340.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 1226.300 2712.070 1340.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2802.470 1340.720 2805.570 1776.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 1776.300 192.070 1890.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 1776.300 372.070 1890.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 1776.300 552.070 1890.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 1776.300 732.070 1890.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 1776.300 2172.070 1890.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 1776.300 2352.070 1890.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 1776.300 2532.070 1890.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 1776.300 2712.070 1890.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2802.470 1890.160 2805.570 2325.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 2326.300 192.070 2940.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 2326.300 372.070 2940.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 2326.300 552.070 2940.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 2326.300 732.070 2940.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 10.640 912.070 2940.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 10.640 1092.070 2940.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 10.640 1272.070 2940.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1448.970 10.640 1452.070 2940.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 10.640 1812.070 2940.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 10.640 1992.070 2940.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 2326.300 2172.070 2940.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 822.470 2940.080 825.570 3375.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.970 10.640 12.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 3376.300 192.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 3376.300 372.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 3376.300 552.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 3376.300 732.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 3376.300 912.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 3376.300 1092.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 3376.300 1272.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1448.970 3376.300 1452.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1628.970 10.640 1632.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 3357.260 1812.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 3357.260 1992.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 3357.260 2172.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 2326.300 2352.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 2326.300 2532.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 2326.300 2712.070 3468.240 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 104.090 2874.080 107.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 284.090 2874.080 287.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 464.090 2874.080 467.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 644.090 2874.080 647.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 98.970 729.390 642.070 732.490 ;
    END
    PORT
      LAYER met5 ;
        RECT 2078.970 729.390 2622.070 732.490 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 824.090 2874.080 827.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 1004.090 2874.080 1007.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 1184.090 2874.080 1187.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 98.970 1278.790 642.070 1281.890 ;
    END
    PORT
      LAYER met5 ;
        RECT 2078.970 1278.790 2622.070 1281.890 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 1364.090 2874.080 1367.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 1544.090 2874.080 1547.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 1724.090 2874.080 1727.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 98.970 1818.790 642.070 1821.890 ;
    END
    PORT
      LAYER met5 ;
        RECT 2078.970 1818.790 2622.070 1821.890 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 1904.090 2874.080 1907.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 2084.090 2874.080 2087.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 2264.090 2874.080 2267.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 2444.090 2874.080 2447.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 2624.090 2874.080 2627.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 2804.090 2874.080 2807.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 2984.090 2874.080 2987.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 3164.090 2874.080 3167.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 3344.090 2874.080 3347.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 98.970 3429.390 1542.070 3432.490 ;
    END
    PORT
      LAYER met5 ;
        RECT 1718.970 3429.390 2082.070 3432.490 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 10.640 102.070 240.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 10.640 282.070 240.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 10.640 462.070 240.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 10.640 642.070 240.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 10.640 2082.070 240.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 10.640 2262.070 240.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 10.640 2442.070 240.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 10.640 2622.070 240.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 12.470 244.560 15.570 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 676.300 102.070 790.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 676.300 282.070 790.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 676.300 462.070 790.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 676.300 642.070 790.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 676.300 2082.070 790.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 676.300 2262.070 790.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 676.300 2442.070 790.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 676.300 2622.070 790.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 12.470 794.000 15.570 1224.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 1226.300 102.070 1340.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 1226.300 282.070 1340.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 1226.300 462.070 1340.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 1226.300 642.070 1340.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 1226.300 2082.070 1340.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 1226.300 2262.070 1340.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 1226.300 2442.070 1340.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 1226.300 2622.070 1340.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 12.470 1343.440 15.570 1773.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 1776.300 102.070 1890.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 1776.300 282.070 1890.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 1776.300 462.070 1890.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 1776.300 642.070 1890.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 1776.300 2082.070 1890.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 1776.300 2262.070 1890.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 1776.300 2442.070 1890.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 1776.300 2622.070 1890.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 12.470 1892.880 15.570 2323.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 2326.300 102.070 2940.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 2326.300 282.070 2940.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 2326.300 462.070 2940.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 2326.300 642.070 2940.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.970 10.640 1002.070 2940.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1178.970 10.640 1182.070 2940.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 10.640 1362.070 2940.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1538.970 10.640 1542.070 2940.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 10.640 1722.070 2940.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 10.640 1902.070 2940.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 2326.300 2082.070 2940.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1632.470 2942.800 1635.570 3356.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 12.470 2942.800 15.570 3373.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 3376.300 102.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 3376.300 282.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 3376.300 462.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 3376.300 642.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.970 10.640 822.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.970 3376.300 1002.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1178.970 3376.300 1182.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 3376.300 1362.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1538.970 3376.300 1542.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 3357.260 1722.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 3357.260 1902.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 3357.260 2082.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 2326.300 2262.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 2326.300 2442.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 2326.300 2622.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2798.970 10.640 2802.070 3468.240 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 1.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 -4.800 8.790 1.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 1.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.670 -4.800 38.230 1.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.470 -4.800 236.030 1.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.950 -4.800 253.510 1.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.890 -4.800 271.450 1.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.370 -4.800 288.930 1.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.850 -4.800 306.410 1.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.330 -4.800 323.890 1.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.810 -4.800 341.370 1.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.290 -4.800 358.850 1.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.770 -4.800 376.330 1.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.250 -4.800 393.810 1.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.670 -4.800 61.230 1.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.730 -4.800 411.290 1.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.210 -4.800 428.770 1.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 -4.800 446.250 1.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.170 -4.800 463.730 1.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.650 -4.800 481.210 1.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.130 -4.800 498.690 1.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.610 -4.800 516.170 1.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.090 -4.800 533.650 1.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.570 -4.800 551.130 1.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.050 -4.800 568.610 1.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.130 -4.800 84.690 1.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.530 -4.800 586.090 1.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.010 -4.800 603.570 1.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.590 -4.800 108.150 1.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.590 -4.800 131.150 1.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.070 -4.800 148.630 1.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.550 -4.800 166.110 1.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.030 -4.800 183.590 1.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.510 -4.800 201.070 1.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.990 -4.800 218.550 1.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 1.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.190 -4.800 43.750 1.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.450 -4.800 242.010 1.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.930 -4.800 259.490 1.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.410 -4.800 276.970 1.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.890 -4.800 294.450 1.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.370 -4.800 311.930 1.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.850 -4.800 329.410 1.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.330 -4.800 346.890 1.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.810 -4.800 364.370 1.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.290 -4.800 381.850 1.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.770 -4.800 399.330 1.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.650 -4.800 67.210 1.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.250 -4.800 416.810 1.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.730 -4.800 434.290 1.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.210 -4.800 451.770 1.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.690 -4.800 469.250 1.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.170 -4.800 486.730 1.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.650 -4.800 504.210 1.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.130 -4.800 521.690 1.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.070 -4.800 539.630 1.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.550 -4.800 557.110 1.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.030 -4.800 574.590 1.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.110 -4.800 90.670 1.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.510 -4.800 592.070 1.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.990 -4.800 609.550 1.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.110 -4.800 113.670 1.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.570 -4.800 137.130 1.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.050 -4.800 154.610 1.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.530 -4.800 172.090 1.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.010 -4.800 189.570 1.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.490 -4.800 207.050 1.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.970 -4.800 224.530 1.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.170 -4.800 49.730 1.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.430 -4.800 247.990 1.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.910 -4.800 265.470 1.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.390 -4.800 282.950 1.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.870 -4.800 300.430 1.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.350 -4.800 317.910 1.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.830 -4.800 335.390 1.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.310 -4.800 352.870 1.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.790 -4.800 370.350 1.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.270 -4.800 387.830 1.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.750 -4.800 405.310 1.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.630 -4.800 73.190 1.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.230 -4.800 422.790 1.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.710 -4.800 440.270 1.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.190 -4.800 457.750 1.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.670 -4.800 475.230 1.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.150 -4.800 492.710 1.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.630 -4.800 510.190 1.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.110 -4.800 527.670 1.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.590 -4.800 545.150 1.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.070 -4.800 562.630 1.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.550 -4.800 580.110 1.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.630 -4.800 96.190 1.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.030 -4.800 597.590 1.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.510 -4.800 615.070 1.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.090 -4.800 119.650 1.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.550 -4.800 143.110 1.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.030 -4.800 160.590 1.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.510 -4.800 178.070 1.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.990 -4.800 195.550 1.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.470 -4.800 213.030 1.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.950 -4.800 230.510 1.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.150 -4.800 55.710 1.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.150 -4.800 78.710 1.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.610 -4.800 102.170 1.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.070 -4.800 125.630 1.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.710 -4.800 26.270 1.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.690 -4.800 32.250 1.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2874.080 3468.085 ;
      LAYER met1 ;
        RECT 2.830 2.420 2877.230 3468.240 ;
      LAYER met2 ;
        RECT 2.860 3478.720 39.230 3479.000 ;
        RECT 40.350 3478.720 118.810 3479.000 ;
        RECT 119.930 3478.720 198.850 3479.000 ;
        RECT 199.970 3478.720 278.890 3479.000 ;
        RECT 280.010 3478.720 358.930 3479.000 ;
        RECT 360.050 3478.720 438.970 3479.000 ;
        RECT 440.090 3478.720 519.010 3479.000 ;
        RECT 520.130 3478.720 599.050 3479.000 ;
        RECT 600.170 3478.720 679.090 3479.000 ;
        RECT 680.210 3478.720 759.130 3479.000 ;
        RECT 760.250 3478.720 839.170 3479.000 ;
        RECT 840.290 3478.720 919.210 3479.000 ;
        RECT 920.330 3478.720 999.250 3479.000 ;
        RECT 1000.370 3478.720 1078.830 3479.000 ;
        RECT 1079.950 3478.720 1158.870 3479.000 ;
        RECT 1159.990 3478.720 1238.910 3479.000 ;
        RECT 1240.030 3478.720 1318.950 3479.000 ;
        RECT 1320.070 3478.720 1398.990 3479.000 ;
        RECT 1400.110 3478.720 1479.030 3479.000 ;
        RECT 1480.150 3478.720 1559.070 3479.000 ;
        RECT 1560.190 3478.720 1639.110 3479.000 ;
        RECT 1640.230 3478.720 1719.150 3479.000 ;
        RECT 1720.270 3478.720 1799.190 3479.000 ;
        RECT 1800.310 3478.720 1879.230 3479.000 ;
        RECT 1880.350 3478.720 1959.270 3479.000 ;
        RECT 1960.390 3478.720 2038.850 3479.000 ;
        RECT 2039.970 3478.720 2118.890 3479.000 ;
        RECT 2120.010 3478.720 2198.930 3479.000 ;
        RECT 2200.050 3478.720 2278.970 3479.000 ;
        RECT 2280.090 3478.720 2359.010 3479.000 ;
        RECT 2360.130 3478.720 2439.050 3479.000 ;
        RECT 2440.170 3478.720 2519.090 3479.000 ;
        RECT 2520.210 3478.720 2599.130 3479.000 ;
        RECT 2600.250 3478.720 2679.170 3479.000 ;
        RECT 2680.290 3478.720 2759.210 3479.000 ;
        RECT 2760.330 3478.720 2839.250 3479.000 ;
        RECT 2840.370 3478.720 2877.200 3479.000 ;
        RECT 2.860 1.280 2877.200 3478.720 ;
        RECT 3.550 0.270 7.950 1.280 ;
        RECT 9.070 0.270 13.930 1.280 ;
        RECT 15.050 0.270 19.910 1.280 ;
        RECT 21.030 0.270 25.430 1.280 ;
        RECT 26.550 0.270 31.410 1.280 ;
        RECT 32.530 0.270 37.390 1.280 ;
        RECT 38.510 0.270 42.910 1.280 ;
        RECT 44.030 0.270 48.890 1.280 ;
        RECT 50.010 0.270 54.870 1.280 ;
        RECT 55.990 0.270 60.390 1.280 ;
        RECT 61.510 0.270 66.370 1.280 ;
        RECT 67.490 0.270 72.350 1.280 ;
        RECT 73.470 0.270 77.870 1.280 ;
        RECT 78.990 0.270 83.850 1.280 ;
        RECT 84.970 0.270 89.830 1.280 ;
        RECT 90.950 0.270 95.350 1.280 ;
        RECT 96.470 0.270 101.330 1.280 ;
        RECT 102.450 0.270 107.310 1.280 ;
        RECT 108.430 0.270 112.830 1.280 ;
        RECT 113.950 0.270 118.810 1.280 ;
        RECT 119.930 0.270 124.790 1.280 ;
        RECT 125.910 0.270 130.310 1.280 ;
        RECT 131.430 0.270 136.290 1.280 ;
        RECT 137.410 0.270 142.270 1.280 ;
        RECT 143.390 0.270 147.790 1.280 ;
        RECT 148.910 0.270 153.770 1.280 ;
        RECT 154.890 0.270 159.750 1.280 ;
        RECT 160.870 0.270 165.270 1.280 ;
        RECT 166.390 0.270 171.250 1.280 ;
        RECT 172.370 0.270 177.230 1.280 ;
        RECT 178.350 0.270 182.750 1.280 ;
        RECT 183.870 0.270 188.730 1.280 ;
        RECT 189.850 0.270 194.710 1.280 ;
        RECT 195.830 0.270 200.230 1.280 ;
        RECT 201.350 0.270 206.210 1.280 ;
        RECT 207.330 0.270 212.190 1.280 ;
        RECT 213.310 0.270 217.710 1.280 ;
        RECT 218.830 0.270 223.690 1.280 ;
        RECT 224.810 0.270 229.670 1.280 ;
        RECT 230.790 0.270 235.190 1.280 ;
        RECT 236.310 0.270 241.170 1.280 ;
        RECT 242.290 0.270 247.150 1.280 ;
        RECT 248.270 0.270 252.670 1.280 ;
        RECT 253.790 0.270 258.650 1.280 ;
        RECT 259.770 0.270 264.630 1.280 ;
        RECT 265.750 0.270 270.610 1.280 ;
        RECT 271.730 0.270 276.130 1.280 ;
        RECT 277.250 0.270 282.110 1.280 ;
        RECT 283.230 0.270 288.090 1.280 ;
        RECT 289.210 0.270 293.610 1.280 ;
        RECT 294.730 0.270 299.590 1.280 ;
        RECT 300.710 0.270 305.570 1.280 ;
        RECT 306.690 0.270 311.090 1.280 ;
        RECT 312.210 0.270 317.070 1.280 ;
        RECT 318.190 0.270 323.050 1.280 ;
        RECT 324.170 0.270 328.570 1.280 ;
        RECT 329.690 0.270 334.550 1.280 ;
        RECT 335.670 0.270 340.530 1.280 ;
        RECT 341.650 0.270 346.050 1.280 ;
        RECT 347.170 0.270 352.030 1.280 ;
        RECT 353.150 0.270 358.010 1.280 ;
        RECT 359.130 0.270 363.530 1.280 ;
        RECT 364.650 0.270 369.510 1.280 ;
        RECT 370.630 0.270 375.490 1.280 ;
        RECT 376.610 0.270 381.010 1.280 ;
        RECT 382.130 0.270 386.990 1.280 ;
        RECT 388.110 0.270 392.970 1.280 ;
        RECT 394.090 0.270 398.490 1.280 ;
        RECT 399.610 0.270 404.470 1.280 ;
        RECT 405.590 0.270 410.450 1.280 ;
        RECT 411.570 0.270 415.970 1.280 ;
        RECT 417.090 0.270 421.950 1.280 ;
        RECT 423.070 0.270 427.930 1.280 ;
        RECT 429.050 0.270 433.450 1.280 ;
        RECT 434.570 0.270 439.430 1.280 ;
        RECT 440.550 0.270 445.410 1.280 ;
        RECT 446.530 0.270 450.930 1.280 ;
        RECT 452.050 0.270 456.910 1.280 ;
        RECT 458.030 0.270 462.890 1.280 ;
        RECT 464.010 0.270 468.410 1.280 ;
        RECT 469.530 0.270 474.390 1.280 ;
        RECT 475.510 0.270 480.370 1.280 ;
        RECT 481.490 0.270 485.890 1.280 ;
        RECT 487.010 0.270 491.870 1.280 ;
        RECT 492.990 0.270 497.850 1.280 ;
        RECT 498.970 0.270 503.370 1.280 ;
        RECT 504.490 0.270 509.350 1.280 ;
        RECT 510.470 0.270 515.330 1.280 ;
        RECT 516.450 0.270 520.850 1.280 ;
        RECT 521.970 0.270 526.830 1.280 ;
        RECT 527.950 0.270 532.810 1.280 ;
        RECT 533.930 0.270 538.790 1.280 ;
        RECT 539.910 0.270 544.310 1.280 ;
        RECT 545.430 0.270 550.290 1.280 ;
        RECT 551.410 0.270 556.270 1.280 ;
        RECT 557.390 0.270 561.790 1.280 ;
        RECT 562.910 0.270 567.770 1.280 ;
        RECT 568.890 0.270 573.750 1.280 ;
        RECT 574.870 0.270 579.270 1.280 ;
        RECT 580.390 0.270 585.250 1.280 ;
        RECT 586.370 0.270 591.230 1.280 ;
        RECT 592.350 0.270 596.750 1.280 ;
        RECT 597.870 0.270 602.730 1.280 ;
        RECT 603.850 0.270 608.710 1.280 ;
        RECT 609.830 0.270 614.230 1.280 ;
        RECT 615.350 0.270 620.210 1.280 ;
        RECT 621.330 0.270 626.190 1.280 ;
        RECT 627.310 0.270 631.710 1.280 ;
        RECT 632.830 0.270 637.690 1.280 ;
        RECT 638.810 0.270 643.670 1.280 ;
        RECT 644.790 0.270 649.190 1.280 ;
        RECT 650.310 0.270 655.170 1.280 ;
        RECT 656.290 0.270 661.150 1.280 ;
        RECT 662.270 0.270 666.670 1.280 ;
        RECT 667.790 0.270 672.650 1.280 ;
        RECT 673.770 0.270 678.630 1.280 ;
        RECT 679.750 0.270 684.150 1.280 ;
        RECT 685.270 0.270 690.130 1.280 ;
        RECT 691.250 0.270 696.110 1.280 ;
        RECT 697.230 0.270 701.630 1.280 ;
        RECT 702.750 0.270 707.610 1.280 ;
        RECT 708.730 0.270 713.590 1.280 ;
        RECT 714.710 0.270 719.110 1.280 ;
        RECT 720.230 0.270 725.090 1.280 ;
        RECT 726.210 0.270 731.070 1.280 ;
        RECT 732.190 0.270 736.590 1.280 ;
        RECT 737.710 0.270 742.570 1.280 ;
        RECT 743.690 0.270 748.550 1.280 ;
        RECT 749.670 0.270 754.070 1.280 ;
        RECT 755.190 0.270 760.050 1.280 ;
        RECT 761.170 0.270 766.030 1.280 ;
        RECT 767.150 0.270 771.550 1.280 ;
        RECT 772.670 0.270 777.530 1.280 ;
        RECT 778.650 0.270 783.510 1.280 ;
        RECT 784.630 0.270 789.490 1.280 ;
        RECT 790.610 0.270 795.010 1.280 ;
        RECT 796.130 0.270 800.990 1.280 ;
        RECT 802.110 0.270 806.970 1.280 ;
        RECT 808.090 0.270 812.490 1.280 ;
        RECT 813.610 0.270 818.470 1.280 ;
        RECT 819.590 0.270 824.450 1.280 ;
        RECT 825.570 0.270 829.970 1.280 ;
        RECT 831.090 0.270 835.950 1.280 ;
        RECT 837.070 0.270 841.930 1.280 ;
        RECT 843.050 0.270 847.450 1.280 ;
        RECT 848.570 0.270 853.430 1.280 ;
        RECT 854.550 0.270 859.410 1.280 ;
        RECT 860.530 0.270 864.930 1.280 ;
        RECT 866.050 0.270 870.910 1.280 ;
        RECT 872.030 0.270 876.890 1.280 ;
        RECT 878.010 0.270 882.410 1.280 ;
        RECT 883.530 0.270 888.390 1.280 ;
        RECT 889.510 0.270 894.370 1.280 ;
        RECT 895.490 0.270 899.890 1.280 ;
        RECT 901.010 0.270 905.870 1.280 ;
        RECT 906.990 0.270 911.850 1.280 ;
        RECT 912.970 0.270 917.370 1.280 ;
        RECT 918.490 0.270 923.350 1.280 ;
        RECT 924.470 0.270 929.330 1.280 ;
        RECT 930.450 0.270 934.850 1.280 ;
        RECT 935.970 0.270 940.830 1.280 ;
        RECT 941.950 0.270 946.810 1.280 ;
        RECT 947.930 0.270 952.330 1.280 ;
        RECT 953.450 0.270 958.310 1.280 ;
        RECT 959.430 0.270 964.290 1.280 ;
        RECT 965.410 0.270 969.810 1.280 ;
        RECT 970.930 0.270 975.790 1.280 ;
        RECT 976.910 0.270 981.770 1.280 ;
        RECT 982.890 0.270 987.290 1.280 ;
        RECT 988.410 0.270 993.270 1.280 ;
        RECT 994.390 0.270 999.250 1.280 ;
        RECT 1000.370 0.270 1004.770 1.280 ;
        RECT 1005.890 0.270 1010.750 1.280 ;
        RECT 1011.870 0.270 1016.730 1.280 ;
        RECT 1017.850 0.270 1022.250 1.280 ;
        RECT 1023.370 0.270 1028.230 1.280 ;
        RECT 1029.350 0.270 1034.210 1.280 ;
        RECT 1035.330 0.270 1039.730 1.280 ;
        RECT 1040.850 0.270 1045.710 1.280 ;
        RECT 1046.830 0.270 1051.690 1.280 ;
        RECT 1052.810 0.270 1057.670 1.280 ;
        RECT 1058.790 0.270 1063.190 1.280 ;
        RECT 1064.310 0.270 1069.170 1.280 ;
        RECT 1070.290 0.270 1075.150 1.280 ;
        RECT 1076.270 0.270 1080.670 1.280 ;
        RECT 1081.790 0.270 1086.650 1.280 ;
        RECT 1087.770 0.270 1092.630 1.280 ;
        RECT 1093.750 0.270 1098.150 1.280 ;
        RECT 1099.270 0.270 1104.130 1.280 ;
        RECT 1105.250 0.270 1110.110 1.280 ;
        RECT 1111.230 0.270 1115.630 1.280 ;
        RECT 1116.750 0.270 1121.610 1.280 ;
        RECT 1122.730 0.270 1127.590 1.280 ;
        RECT 1128.710 0.270 1133.110 1.280 ;
        RECT 1134.230 0.270 1139.090 1.280 ;
        RECT 1140.210 0.270 1145.070 1.280 ;
        RECT 1146.190 0.270 1150.590 1.280 ;
        RECT 1151.710 0.270 1156.570 1.280 ;
        RECT 1157.690 0.270 1162.550 1.280 ;
        RECT 1163.670 0.270 1168.070 1.280 ;
        RECT 1169.190 0.270 1174.050 1.280 ;
        RECT 1175.170 0.270 1180.030 1.280 ;
        RECT 1181.150 0.270 1185.550 1.280 ;
        RECT 1186.670 0.270 1191.530 1.280 ;
        RECT 1192.650 0.270 1197.510 1.280 ;
        RECT 1198.630 0.270 1203.030 1.280 ;
        RECT 1204.150 0.270 1209.010 1.280 ;
        RECT 1210.130 0.270 1214.990 1.280 ;
        RECT 1216.110 0.270 1220.510 1.280 ;
        RECT 1221.630 0.270 1226.490 1.280 ;
        RECT 1227.610 0.270 1232.470 1.280 ;
        RECT 1233.590 0.270 1237.990 1.280 ;
        RECT 1239.110 0.270 1243.970 1.280 ;
        RECT 1245.090 0.270 1249.950 1.280 ;
        RECT 1251.070 0.270 1255.470 1.280 ;
        RECT 1256.590 0.270 1261.450 1.280 ;
        RECT 1262.570 0.270 1267.430 1.280 ;
        RECT 1268.550 0.270 1272.950 1.280 ;
        RECT 1274.070 0.270 1278.930 1.280 ;
        RECT 1280.050 0.270 1284.910 1.280 ;
        RECT 1286.030 0.270 1290.430 1.280 ;
        RECT 1291.550 0.270 1296.410 1.280 ;
        RECT 1297.530 0.270 1302.390 1.280 ;
        RECT 1303.510 0.270 1307.910 1.280 ;
        RECT 1309.030 0.270 1313.890 1.280 ;
        RECT 1315.010 0.270 1319.870 1.280 ;
        RECT 1320.990 0.270 1325.850 1.280 ;
        RECT 1326.970 0.270 1331.370 1.280 ;
        RECT 1332.490 0.270 1337.350 1.280 ;
        RECT 1338.470 0.270 1343.330 1.280 ;
        RECT 1344.450 0.270 1348.850 1.280 ;
        RECT 1349.970 0.270 1354.830 1.280 ;
        RECT 1355.950 0.270 1360.810 1.280 ;
        RECT 1361.930 0.270 1366.330 1.280 ;
        RECT 1367.450 0.270 1372.310 1.280 ;
        RECT 1373.430 0.270 1378.290 1.280 ;
        RECT 1379.410 0.270 1383.810 1.280 ;
        RECT 1384.930 0.270 1389.790 1.280 ;
        RECT 1390.910 0.270 1395.770 1.280 ;
        RECT 1396.890 0.270 1401.290 1.280 ;
        RECT 1402.410 0.270 1407.270 1.280 ;
        RECT 1408.390 0.270 1413.250 1.280 ;
        RECT 1414.370 0.270 1418.770 1.280 ;
        RECT 1419.890 0.270 1424.750 1.280 ;
        RECT 1425.870 0.270 1430.730 1.280 ;
        RECT 1431.850 0.270 1436.250 1.280 ;
        RECT 1437.370 0.270 1442.230 1.280 ;
        RECT 1443.350 0.270 1448.210 1.280 ;
        RECT 1449.330 0.270 1453.730 1.280 ;
        RECT 1454.850 0.270 1459.710 1.280 ;
        RECT 1460.830 0.270 1465.690 1.280 ;
        RECT 1466.810 0.270 1471.210 1.280 ;
        RECT 1472.330 0.270 1477.190 1.280 ;
        RECT 1478.310 0.270 1483.170 1.280 ;
        RECT 1484.290 0.270 1488.690 1.280 ;
        RECT 1489.810 0.270 1494.670 1.280 ;
        RECT 1495.790 0.270 1500.650 1.280 ;
        RECT 1501.770 0.270 1506.170 1.280 ;
        RECT 1507.290 0.270 1512.150 1.280 ;
        RECT 1513.270 0.270 1518.130 1.280 ;
        RECT 1519.250 0.270 1523.650 1.280 ;
        RECT 1524.770 0.270 1529.630 1.280 ;
        RECT 1530.750 0.270 1535.610 1.280 ;
        RECT 1536.730 0.270 1541.130 1.280 ;
        RECT 1542.250 0.270 1547.110 1.280 ;
        RECT 1548.230 0.270 1553.090 1.280 ;
        RECT 1554.210 0.270 1558.610 1.280 ;
        RECT 1559.730 0.270 1564.590 1.280 ;
        RECT 1565.710 0.270 1570.570 1.280 ;
        RECT 1571.690 0.270 1576.550 1.280 ;
        RECT 1577.670 0.270 1582.070 1.280 ;
        RECT 1583.190 0.270 1588.050 1.280 ;
        RECT 1589.170 0.270 1594.030 1.280 ;
        RECT 1595.150 0.270 1599.550 1.280 ;
        RECT 1600.670 0.270 1605.530 1.280 ;
        RECT 1606.650 0.270 1611.510 1.280 ;
        RECT 1612.630 0.270 1617.030 1.280 ;
        RECT 1618.150 0.270 1623.010 1.280 ;
        RECT 1624.130 0.270 1628.990 1.280 ;
        RECT 1630.110 0.270 1634.510 1.280 ;
        RECT 1635.630 0.270 1640.490 1.280 ;
        RECT 1641.610 0.270 1646.470 1.280 ;
        RECT 1647.590 0.270 1651.990 1.280 ;
        RECT 1653.110 0.270 1657.970 1.280 ;
        RECT 1659.090 0.270 1663.950 1.280 ;
        RECT 1665.070 0.270 1669.470 1.280 ;
        RECT 1670.590 0.270 1675.450 1.280 ;
        RECT 1676.570 0.270 1681.430 1.280 ;
        RECT 1682.550 0.270 1686.950 1.280 ;
        RECT 1688.070 0.270 1692.930 1.280 ;
        RECT 1694.050 0.270 1698.910 1.280 ;
        RECT 1700.030 0.270 1704.430 1.280 ;
        RECT 1705.550 0.270 1710.410 1.280 ;
        RECT 1711.530 0.270 1716.390 1.280 ;
        RECT 1717.510 0.270 1721.910 1.280 ;
        RECT 1723.030 0.270 1727.890 1.280 ;
        RECT 1729.010 0.270 1733.870 1.280 ;
        RECT 1734.990 0.270 1739.390 1.280 ;
        RECT 1740.510 0.270 1745.370 1.280 ;
        RECT 1746.490 0.270 1751.350 1.280 ;
        RECT 1752.470 0.270 1756.870 1.280 ;
        RECT 1757.990 0.270 1762.850 1.280 ;
        RECT 1763.970 0.270 1768.830 1.280 ;
        RECT 1769.950 0.270 1774.350 1.280 ;
        RECT 1775.470 0.270 1780.330 1.280 ;
        RECT 1781.450 0.270 1786.310 1.280 ;
        RECT 1787.430 0.270 1791.830 1.280 ;
        RECT 1792.950 0.270 1797.810 1.280 ;
        RECT 1798.930 0.270 1803.790 1.280 ;
        RECT 1804.910 0.270 1809.310 1.280 ;
        RECT 1810.430 0.270 1815.290 1.280 ;
        RECT 1816.410 0.270 1821.270 1.280 ;
        RECT 1822.390 0.270 1826.790 1.280 ;
        RECT 1827.910 0.270 1832.770 1.280 ;
        RECT 1833.890 0.270 1838.750 1.280 ;
        RECT 1839.870 0.270 1844.730 1.280 ;
        RECT 1845.850 0.270 1850.250 1.280 ;
        RECT 1851.370 0.270 1856.230 1.280 ;
        RECT 1857.350 0.270 1862.210 1.280 ;
        RECT 1863.330 0.270 1867.730 1.280 ;
        RECT 1868.850 0.270 1873.710 1.280 ;
        RECT 1874.830 0.270 1879.690 1.280 ;
        RECT 1880.810 0.270 1885.210 1.280 ;
        RECT 1886.330 0.270 1891.190 1.280 ;
        RECT 1892.310 0.270 1897.170 1.280 ;
        RECT 1898.290 0.270 1902.690 1.280 ;
        RECT 1903.810 0.270 1908.670 1.280 ;
        RECT 1909.790 0.270 1914.650 1.280 ;
        RECT 1915.770 0.270 1920.170 1.280 ;
        RECT 1921.290 0.270 1926.150 1.280 ;
        RECT 1927.270 0.270 1932.130 1.280 ;
        RECT 1933.250 0.270 1937.650 1.280 ;
        RECT 1938.770 0.270 1943.630 1.280 ;
        RECT 1944.750 0.270 1949.610 1.280 ;
        RECT 1950.730 0.270 1955.130 1.280 ;
        RECT 1956.250 0.270 1961.110 1.280 ;
        RECT 1962.230 0.270 1967.090 1.280 ;
        RECT 1968.210 0.270 1972.610 1.280 ;
        RECT 1973.730 0.270 1978.590 1.280 ;
        RECT 1979.710 0.270 1984.570 1.280 ;
        RECT 1985.690 0.270 1990.090 1.280 ;
        RECT 1991.210 0.270 1996.070 1.280 ;
        RECT 1997.190 0.270 2002.050 1.280 ;
        RECT 2003.170 0.270 2007.570 1.280 ;
        RECT 2008.690 0.270 2013.550 1.280 ;
        RECT 2014.670 0.270 2019.530 1.280 ;
        RECT 2020.650 0.270 2025.050 1.280 ;
        RECT 2026.170 0.270 2031.030 1.280 ;
        RECT 2032.150 0.270 2037.010 1.280 ;
        RECT 2038.130 0.270 2042.530 1.280 ;
        RECT 2043.650 0.270 2048.510 1.280 ;
        RECT 2049.630 0.270 2054.490 1.280 ;
        RECT 2055.610 0.270 2060.010 1.280 ;
        RECT 2061.130 0.270 2065.990 1.280 ;
        RECT 2067.110 0.270 2071.970 1.280 ;
        RECT 2073.090 0.270 2077.490 1.280 ;
        RECT 2078.610 0.270 2083.470 1.280 ;
        RECT 2084.590 0.270 2089.450 1.280 ;
        RECT 2090.570 0.270 2094.970 1.280 ;
        RECT 2096.090 0.270 2100.950 1.280 ;
        RECT 2102.070 0.270 2106.930 1.280 ;
        RECT 2108.050 0.270 2112.910 1.280 ;
        RECT 2114.030 0.270 2118.430 1.280 ;
        RECT 2119.550 0.270 2124.410 1.280 ;
        RECT 2125.530 0.270 2130.390 1.280 ;
        RECT 2131.510 0.270 2135.910 1.280 ;
        RECT 2137.030 0.270 2141.890 1.280 ;
        RECT 2143.010 0.270 2147.870 1.280 ;
        RECT 2148.990 0.270 2153.390 1.280 ;
        RECT 2154.510 0.270 2159.370 1.280 ;
        RECT 2160.490 0.270 2165.350 1.280 ;
        RECT 2166.470 0.270 2170.870 1.280 ;
        RECT 2171.990 0.270 2176.850 1.280 ;
        RECT 2177.970 0.270 2182.830 1.280 ;
        RECT 2183.950 0.270 2188.350 1.280 ;
        RECT 2189.470 0.270 2194.330 1.280 ;
        RECT 2195.450 0.270 2200.310 1.280 ;
        RECT 2201.430 0.270 2205.830 1.280 ;
        RECT 2206.950 0.270 2211.810 1.280 ;
        RECT 2212.930 0.270 2217.790 1.280 ;
        RECT 2218.910 0.270 2223.310 1.280 ;
        RECT 2224.430 0.270 2229.290 1.280 ;
        RECT 2230.410 0.270 2235.270 1.280 ;
        RECT 2236.390 0.270 2240.790 1.280 ;
        RECT 2241.910 0.270 2246.770 1.280 ;
        RECT 2247.890 0.270 2252.750 1.280 ;
        RECT 2253.870 0.270 2258.270 1.280 ;
        RECT 2259.390 0.270 2264.250 1.280 ;
        RECT 2265.370 0.270 2270.230 1.280 ;
        RECT 2271.350 0.270 2275.750 1.280 ;
        RECT 2276.870 0.270 2281.730 1.280 ;
        RECT 2282.850 0.270 2287.710 1.280 ;
        RECT 2288.830 0.270 2293.230 1.280 ;
        RECT 2294.350 0.270 2299.210 1.280 ;
        RECT 2300.330 0.270 2305.190 1.280 ;
        RECT 2306.310 0.270 2310.710 1.280 ;
        RECT 2311.830 0.270 2316.690 1.280 ;
        RECT 2317.810 0.270 2322.670 1.280 ;
        RECT 2323.790 0.270 2328.190 1.280 ;
        RECT 2329.310 0.270 2334.170 1.280 ;
        RECT 2335.290 0.270 2340.150 1.280 ;
        RECT 2341.270 0.270 2345.670 1.280 ;
        RECT 2346.790 0.270 2351.650 1.280 ;
        RECT 2352.770 0.270 2357.630 1.280 ;
        RECT 2358.750 0.270 2363.610 1.280 ;
        RECT 2364.730 0.270 2369.130 1.280 ;
        RECT 2370.250 0.270 2375.110 1.280 ;
        RECT 2376.230 0.270 2381.090 1.280 ;
        RECT 2382.210 0.270 2386.610 1.280 ;
        RECT 2387.730 0.270 2392.590 1.280 ;
        RECT 2393.710 0.270 2398.570 1.280 ;
        RECT 2399.690 0.270 2404.090 1.280 ;
        RECT 2405.210 0.270 2410.070 1.280 ;
        RECT 2411.190 0.270 2416.050 1.280 ;
        RECT 2417.170 0.270 2421.570 1.280 ;
        RECT 2422.690 0.270 2427.550 1.280 ;
        RECT 2428.670 0.270 2433.530 1.280 ;
        RECT 2434.650 0.270 2439.050 1.280 ;
        RECT 2440.170 0.270 2445.030 1.280 ;
        RECT 2446.150 0.270 2451.010 1.280 ;
        RECT 2452.130 0.270 2456.530 1.280 ;
        RECT 2457.650 0.270 2462.510 1.280 ;
        RECT 2463.630 0.270 2468.490 1.280 ;
        RECT 2469.610 0.270 2474.010 1.280 ;
        RECT 2475.130 0.270 2479.990 1.280 ;
        RECT 2481.110 0.270 2485.970 1.280 ;
        RECT 2487.090 0.270 2491.490 1.280 ;
        RECT 2492.610 0.270 2497.470 1.280 ;
        RECT 2498.590 0.270 2503.450 1.280 ;
        RECT 2504.570 0.270 2508.970 1.280 ;
        RECT 2510.090 0.270 2514.950 1.280 ;
        RECT 2516.070 0.270 2520.930 1.280 ;
        RECT 2522.050 0.270 2526.450 1.280 ;
        RECT 2527.570 0.270 2532.430 1.280 ;
        RECT 2533.550 0.270 2538.410 1.280 ;
        RECT 2539.530 0.270 2543.930 1.280 ;
        RECT 2545.050 0.270 2549.910 1.280 ;
        RECT 2551.030 0.270 2555.890 1.280 ;
        RECT 2557.010 0.270 2561.410 1.280 ;
        RECT 2562.530 0.270 2567.390 1.280 ;
        RECT 2568.510 0.270 2573.370 1.280 ;
        RECT 2574.490 0.270 2578.890 1.280 ;
        RECT 2580.010 0.270 2584.870 1.280 ;
        RECT 2585.990 0.270 2590.850 1.280 ;
        RECT 2591.970 0.270 2596.370 1.280 ;
        RECT 2597.490 0.270 2602.350 1.280 ;
        RECT 2603.470 0.270 2608.330 1.280 ;
        RECT 2609.450 0.270 2613.850 1.280 ;
        RECT 2614.970 0.270 2619.830 1.280 ;
        RECT 2620.950 0.270 2625.810 1.280 ;
        RECT 2626.930 0.270 2631.790 1.280 ;
        RECT 2632.910 0.270 2637.310 1.280 ;
        RECT 2638.430 0.270 2643.290 1.280 ;
        RECT 2644.410 0.270 2649.270 1.280 ;
        RECT 2650.390 0.270 2654.790 1.280 ;
        RECT 2655.910 0.270 2660.770 1.280 ;
        RECT 2661.890 0.270 2666.750 1.280 ;
        RECT 2667.870 0.270 2672.270 1.280 ;
        RECT 2673.390 0.270 2678.250 1.280 ;
        RECT 2679.370 0.270 2684.230 1.280 ;
        RECT 2685.350 0.270 2689.750 1.280 ;
        RECT 2690.870 0.270 2695.730 1.280 ;
        RECT 2696.850 0.270 2701.710 1.280 ;
        RECT 2702.830 0.270 2707.230 1.280 ;
        RECT 2708.350 0.270 2713.210 1.280 ;
        RECT 2714.330 0.270 2719.190 1.280 ;
        RECT 2720.310 0.270 2724.710 1.280 ;
        RECT 2725.830 0.270 2730.690 1.280 ;
        RECT 2731.810 0.270 2736.670 1.280 ;
        RECT 2737.790 0.270 2742.190 1.280 ;
        RECT 2743.310 0.270 2748.170 1.280 ;
        RECT 2749.290 0.270 2754.150 1.280 ;
        RECT 2755.270 0.270 2759.670 1.280 ;
        RECT 2760.790 0.270 2765.650 1.280 ;
        RECT 2766.770 0.270 2771.630 1.280 ;
        RECT 2772.750 0.270 2777.150 1.280 ;
        RECT 2778.270 0.270 2783.130 1.280 ;
        RECT 2784.250 0.270 2789.110 1.280 ;
        RECT 2790.230 0.270 2794.630 1.280 ;
        RECT 2795.750 0.270 2800.610 1.280 ;
        RECT 2801.730 0.270 2806.590 1.280 ;
        RECT 2807.710 0.270 2812.110 1.280 ;
        RECT 2813.230 0.270 2818.090 1.280 ;
        RECT 2819.210 0.270 2824.070 1.280 ;
        RECT 2825.190 0.270 2829.590 1.280 ;
        RECT 2830.710 0.270 2835.570 1.280 ;
        RECT 2836.690 0.270 2841.550 1.280 ;
        RECT 2842.670 0.270 2847.070 1.280 ;
        RECT 2848.190 0.270 2853.050 1.280 ;
        RECT 2854.170 0.270 2859.030 1.280 ;
        RECT 2860.150 0.270 2864.550 1.280 ;
        RECT 2865.670 0.270 2870.530 1.280 ;
        RECT 2871.650 0.270 2876.510 1.280 ;
      LAYER met3 ;
        RECT 1.000 3448.940 2879.000 3468.165 ;
        RECT 1.400 3448.260 2879.000 3448.940 ;
        RECT 1.400 3446.940 2878.600 3448.260 ;
        RECT 1.000 3446.260 2878.600 3446.940 ;
        RECT 1.000 3384.340 2879.000 3446.260 ;
        RECT 1.400 3382.340 2879.000 3384.340 ;
        RECT 1.000 3382.300 2879.000 3382.340 ;
        RECT 1.000 3380.300 2878.600 3382.300 ;
        RECT 1.000 3319.740 2879.000 3380.300 ;
        RECT 1.400 3317.740 2879.000 3319.740 ;
        RECT 1.000 3317.020 2879.000 3317.740 ;
        RECT 1.000 3315.020 2878.600 3317.020 ;
        RECT 1.000 3255.140 2879.000 3315.020 ;
        RECT 1.400 3253.140 2879.000 3255.140 ;
        RECT 1.000 3251.060 2879.000 3253.140 ;
        RECT 1.000 3249.060 2878.600 3251.060 ;
        RECT 1.000 3191.220 2879.000 3249.060 ;
        RECT 1.400 3189.220 2879.000 3191.220 ;
        RECT 1.000 3185.780 2879.000 3189.220 ;
        RECT 1.000 3183.780 2878.600 3185.780 ;
        RECT 1.000 3126.620 2879.000 3183.780 ;
        RECT 1.400 3124.620 2879.000 3126.620 ;
        RECT 1.000 3119.820 2879.000 3124.620 ;
        RECT 1.000 3117.820 2878.600 3119.820 ;
        RECT 1.000 3062.020 2879.000 3117.820 ;
        RECT 1.400 3060.020 2879.000 3062.020 ;
        RECT 1.000 3054.540 2879.000 3060.020 ;
        RECT 1.000 3052.540 2878.600 3054.540 ;
        RECT 1.000 2997.420 2879.000 3052.540 ;
        RECT 1.400 2995.420 2879.000 2997.420 ;
        RECT 1.000 2988.580 2879.000 2995.420 ;
        RECT 1.000 2986.580 2878.600 2988.580 ;
        RECT 1.000 2933.500 2879.000 2986.580 ;
        RECT 1.400 2931.500 2879.000 2933.500 ;
        RECT 1.000 2922.620 2879.000 2931.500 ;
        RECT 1.000 2920.620 2878.600 2922.620 ;
        RECT 1.000 2868.900 2879.000 2920.620 ;
        RECT 1.400 2866.900 2879.000 2868.900 ;
        RECT 1.000 2857.340 2879.000 2866.900 ;
        RECT 1.000 2855.340 2878.600 2857.340 ;
        RECT 1.000 2804.300 2879.000 2855.340 ;
        RECT 1.400 2802.300 2879.000 2804.300 ;
        RECT 1.000 2791.380 2879.000 2802.300 ;
        RECT 1.000 2789.380 2878.600 2791.380 ;
        RECT 1.000 2739.700 2879.000 2789.380 ;
        RECT 1.400 2737.700 2879.000 2739.700 ;
        RECT 1.000 2726.100 2879.000 2737.700 ;
        RECT 1.000 2724.100 2878.600 2726.100 ;
        RECT 1.000 2675.100 2879.000 2724.100 ;
        RECT 1.400 2673.100 2879.000 2675.100 ;
        RECT 1.000 2660.140 2879.000 2673.100 ;
        RECT 1.000 2658.140 2878.600 2660.140 ;
        RECT 1.000 2611.180 2879.000 2658.140 ;
        RECT 1.400 2609.180 2879.000 2611.180 ;
        RECT 1.000 2594.860 2879.000 2609.180 ;
        RECT 1.000 2592.860 2878.600 2594.860 ;
        RECT 1.000 2546.580 2879.000 2592.860 ;
        RECT 1.400 2544.580 2879.000 2546.580 ;
        RECT 1.000 2528.900 2879.000 2544.580 ;
        RECT 1.000 2526.900 2878.600 2528.900 ;
        RECT 1.000 2481.980 2879.000 2526.900 ;
        RECT 1.400 2479.980 2879.000 2481.980 ;
        RECT 1.000 2462.940 2879.000 2479.980 ;
        RECT 1.000 2460.940 2878.600 2462.940 ;
        RECT 1.000 2417.380 2879.000 2460.940 ;
        RECT 1.400 2415.380 2879.000 2417.380 ;
        RECT 1.000 2397.660 2879.000 2415.380 ;
        RECT 1.000 2395.660 2878.600 2397.660 ;
        RECT 1.000 2353.460 2879.000 2395.660 ;
        RECT 1.400 2351.460 2879.000 2353.460 ;
        RECT 1.000 2331.700 2879.000 2351.460 ;
        RECT 1.000 2329.700 2878.600 2331.700 ;
        RECT 1.000 2288.860 2879.000 2329.700 ;
        RECT 1.400 2286.860 2879.000 2288.860 ;
        RECT 1.000 2266.420 2879.000 2286.860 ;
        RECT 1.000 2264.420 2878.600 2266.420 ;
        RECT 1.000 2224.260 2879.000 2264.420 ;
        RECT 1.400 2222.260 2879.000 2224.260 ;
        RECT 1.000 2200.460 2879.000 2222.260 ;
        RECT 1.000 2198.460 2878.600 2200.460 ;
        RECT 1.000 2159.660 2879.000 2198.460 ;
        RECT 1.400 2157.660 2879.000 2159.660 ;
        RECT 1.000 2135.180 2879.000 2157.660 ;
        RECT 1.000 2133.180 2878.600 2135.180 ;
        RECT 1.000 2095.060 2879.000 2133.180 ;
        RECT 1.400 2093.060 2879.000 2095.060 ;
        RECT 1.000 2069.220 2879.000 2093.060 ;
        RECT 1.000 2067.220 2878.600 2069.220 ;
        RECT 1.000 2031.140 2879.000 2067.220 ;
        RECT 1.400 2029.140 2879.000 2031.140 ;
        RECT 1.000 2003.260 2879.000 2029.140 ;
        RECT 1.000 2001.260 2878.600 2003.260 ;
        RECT 1.000 1966.540 2879.000 2001.260 ;
        RECT 1.400 1964.540 2879.000 1966.540 ;
        RECT 1.000 1937.980 2879.000 1964.540 ;
        RECT 1.000 1935.980 2878.600 1937.980 ;
        RECT 1.000 1901.940 2879.000 1935.980 ;
        RECT 1.400 1899.940 2879.000 1901.940 ;
        RECT 1.000 1872.020 2879.000 1899.940 ;
        RECT 1.000 1870.020 2878.600 1872.020 ;
        RECT 1.000 1837.340 2879.000 1870.020 ;
        RECT 1.400 1835.340 2879.000 1837.340 ;
        RECT 1.000 1806.740 2879.000 1835.340 ;
        RECT 1.000 1804.740 2878.600 1806.740 ;
        RECT 1.000 1773.420 2879.000 1804.740 ;
        RECT 1.400 1771.420 2879.000 1773.420 ;
        RECT 1.000 1740.780 2879.000 1771.420 ;
        RECT 1.000 1738.780 2878.600 1740.780 ;
        RECT 1.000 1708.820 2879.000 1738.780 ;
        RECT 1.400 1706.820 2879.000 1708.820 ;
        RECT 1.000 1675.500 2879.000 1706.820 ;
        RECT 1.000 1673.500 2878.600 1675.500 ;
        RECT 1.000 1644.220 2879.000 1673.500 ;
        RECT 1.400 1642.220 2879.000 1644.220 ;
        RECT 1.000 1609.540 2879.000 1642.220 ;
        RECT 1.000 1607.540 2878.600 1609.540 ;
        RECT 1.000 1579.620 2879.000 1607.540 ;
        RECT 1.400 1577.620 2879.000 1579.620 ;
        RECT 1.000 1544.260 2879.000 1577.620 ;
        RECT 1.000 1542.260 2878.600 1544.260 ;
        RECT 1.000 1515.020 2879.000 1542.260 ;
        RECT 1.400 1513.020 2879.000 1515.020 ;
        RECT 1.000 1478.300 2879.000 1513.020 ;
        RECT 1.000 1476.300 2878.600 1478.300 ;
        RECT 1.000 1451.100 2879.000 1476.300 ;
        RECT 1.400 1449.100 2879.000 1451.100 ;
        RECT 1.000 1412.340 2879.000 1449.100 ;
        RECT 1.000 1410.340 2878.600 1412.340 ;
        RECT 1.000 1386.500 2879.000 1410.340 ;
        RECT 1.400 1384.500 2879.000 1386.500 ;
        RECT 1.000 1347.060 2879.000 1384.500 ;
        RECT 1.000 1345.060 2878.600 1347.060 ;
        RECT 1.000 1321.900 2879.000 1345.060 ;
        RECT 1.400 1319.900 2879.000 1321.900 ;
        RECT 1.000 1281.100 2879.000 1319.900 ;
        RECT 1.000 1279.100 2878.600 1281.100 ;
        RECT 1.000 1257.300 2879.000 1279.100 ;
        RECT 1.400 1255.300 2879.000 1257.300 ;
        RECT 1.000 1215.820 2879.000 1255.300 ;
        RECT 1.000 1213.820 2878.600 1215.820 ;
        RECT 1.000 1193.380 2879.000 1213.820 ;
        RECT 1.400 1191.380 2879.000 1193.380 ;
        RECT 1.000 1149.860 2879.000 1191.380 ;
        RECT 1.000 1147.860 2878.600 1149.860 ;
        RECT 1.000 1128.780 2879.000 1147.860 ;
        RECT 1.400 1126.780 2879.000 1128.780 ;
        RECT 1.000 1084.580 2879.000 1126.780 ;
        RECT 1.000 1082.580 2878.600 1084.580 ;
        RECT 1.000 1064.180 2879.000 1082.580 ;
        RECT 1.400 1062.180 2879.000 1064.180 ;
        RECT 1.000 1018.620 2879.000 1062.180 ;
        RECT 1.000 1016.620 2878.600 1018.620 ;
        RECT 1.000 999.580 2879.000 1016.620 ;
        RECT 1.400 997.580 2879.000 999.580 ;
        RECT 1.000 952.660 2879.000 997.580 ;
        RECT 1.000 950.660 2878.600 952.660 ;
        RECT 1.000 934.980 2879.000 950.660 ;
        RECT 1.400 932.980 2879.000 934.980 ;
        RECT 1.000 887.380 2879.000 932.980 ;
        RECT 1.000 885.380 2878.600 887.380 ;
        RECT 1.000 871.060 2879.000 885.380 ;
        RECT 1.400 869.060 2879.000 871.060 ;
        RECT 1.000 821.420 2879.000 869.060 ;
        RECT 1.000 819.420 2878.600 821.420 ;
        RECT 1.000 806.460 2879.000 819.420 ;
        RECT 1.400 804.460 2879.000 806.460 ;
        RECT 1.000 756.140 2879.000 804.460 ;
        RECT 1.000 754.140 2878.600 756.140 ;
        RECT 1.000 741.860 2879.000 754.140 ;
        RECT 1.400 739.860 2879.000 741.860 ;
        RECT 1.000 690.180 2879.000 739.860 ;
        RECT 1.000 688.180 2878.600 690.180 ;
        RECT 1.000 677.260 2879.000 688.180 ;
        RECT 1.400 675.260 2879.000 677.260 ;
        RECT 1.000 624.900 2879.000 675.260 ;
        RECT 1.000 622.900 2878.600 624.900 ;
        RECT 1.000 613.340 2879.000 622.900 ;
        RECT 1.400 611.340 2879.000 613.340 ;
        RECT 1.000 558.940 2879.000 611.340 ;
        RECT 1.000 556.940 2878.600 558.940 ;
        RECT 1.000 548.740 2879.000 556.940 ;
        RECT 1.400 546.740 2879.000 548.740 ;
        RECT 1.000 492.980 2879.000 546.740 ;
        RECT 1.000 490.980 2878.600 492.980 ;
        RECT 1.000 484.140 2879.000 490.980 ;
        RECT 1.400 482.140 2879.000 484.140 ;
        RECT 1.000 427.700 2879.000 482.140 ;
        RECT 1.000 425.700 2878.600 427.700 ;
        RECT 1.000 419.540 2879.000 425.700 ;
        RECT 1.400 417.540 2879.000 419.540 ;
        RECT 1.000 361.740 2879.000 417.540 ;
        RECT 1.000 359.740 2878.600 361.740 ;
        RECT 1.000 354.940 2879.000 359.740 ;
        RECT 1.400 352.940 2879.000 354.940 ;
        RECT 1.000 296.460 2879.000 352.940 ;
        RECT 1.000 294.460 2878.600 296.460 ;
        RECT 1.000 291.020 2879.000 294.460 ;
        RECT 1.400 289.020 2879.000 291.020 ;
        RECT 1.000 230.500 2879.000 289.020 ;
        RECT 1.000 228.500 2878.600 230.500 ;
        RECT 1.000 226.420 2879.000 228.500 ;
        RECT 1.400 224.420 2879.000 226.420 ;
        RECT 1.000 165.220 2879.000 224.420 ;
        RECT 1.000 163.220 2878.600 165.220 ;
        RECT 1.000 161.820 2879.000 163.220 ;
        RECT 1.400 159.820 2879.000 161.820 ;
        RECT 1.000 99.260 2879.000 159.820 ;
        RECT 1.000 97.260 2878.600 99.260 ;
        RECT 1.000 97.220 2879.000 97.260 ;
        RECT 1.400 95.220 2879.000 97.220 ;
        RECT 1.000 33.980 2879.000 95.220 ;
        RECT 1.000 33.300 2878.600 33.980 ;
        RECT 1.400 31.980 2878.600 33.300 ;
        RECT 1.400 31.300 2879.000 31.980 ;
        RECT 1.000 2.895 2879.000 31.300 ;
      LAYER met4 ;
        RECT 7.230 10.240 8.570 3467.145 ;
        RECT 12.470 3375.900 98.570 3467.145 ;
        RECT 102.470 3375.900 188.570 3467.145 ;
        RECT 192.470 3375.900 278.570 3467.145 ;
        RECT 282.470 3375.900 368.570 3467.145 ;
        RECT 372.470 3375.900 458.570 3467.145 ;
        RECT 462.470 3375.900 548.570 3467.145 ;
        RECT 552.470 3375.900 638.570 3467.145 ;
        RECT 642.470 3375.900 728.570 3467.145 ;
        RECT 732.470 3375.900 818.570 3467.145 ;
        RECT 822.470 3376.160 908.570 3467.145 ;
        RECT 12.470 3373.440 818.570 3375.900 ;
        RECT 15.970 2942.400 818.570 3373.440 ;
        RECT 12.470 2940.640 818.570 2942.400 ;
        RECT 12.470 2325.900 98.570 2940.640 ;
        RECT 102.470 2325.900 188.570 2940.640 ;
        RECT 192.470 2325.900 278.570 2940.640 ;
        RECT 282.470 2325.900 368.570 2940.640 ;
        RECT 372.470 2325.900 458.570 2940.640 ;
        RECT 462.470 2325.900 548.570 2940.640 ;
        RECT 552.470 2325.900 638.570 2940.640 ;
        RECT 642.470 2325.900 728.570 2940.640 ;
        RECT 732.470 2325.900 818.570 2940.640 ;
        RECT 825.970 3375.900 908.570 3376.160 ;
        RECT 912.470 3375.900 998.570 3467.145 ;
        RECT 1002.470 3375.900 1088.570 3467.145 ;
        RECT 1092.470 3375.900 1178.570 3467.145 ;
        RECT 1182.470 3375.900 1268.570 3467.145 ;
        RECT 1272.470 3375.900 1358.570 3467.145 ;
        RECT 1362.470 3375.900 1448.570 3467.145 ;
        RECT 1452.470 3375.900 1538.570 3467.145 ;
        RECT 1542.470 3375.900 1628.570 3467.145 ;
        RECT 825.970 2940.640 1628.570 3375.900 ;
        RECT 1632.470 3357.120 1718.570 3467.145 ;
        RECT 1635.970 3356.860 1718.570 3357.120 ;
        RECT 1722.470 3356.860 1808.570 3467.145 ;
        RECT 1812.470 3356.860 1898.570 3467.145 ;
        RECT 1902.470 3356.860 1988.570 3467.145 ;
        RECT 1992.470 3356.860 2078.570 3467.145 ;
        RECT 2082.470 3356.860 2168.570 3467.145 ;
        RECT 2172.470 3356.860 2258.570 3467.145 ;
        RECT 1635.970 2942.400 2258.570 3356.860 ;
        RECT 825.970 2939.680 908.570 2940.640 ;
        RECT 12.470 2323.520 818.570 2325.900 ;
        RECT 15.970 1892.480 818.570 2323.520 ;
        RECT 12.470 1890.640 818.570 1892.480 ;
        RECT 12.470 1775.900 98.570 1890.640 ;
        RECT 102.470 1775.900 188.570 1890.640 ;
        RECT 192.470 1775.900 278.570 1890.640 ;
        RECT 282.470 1775.900 368.570 1890.640 ;
        RECT 372.470 1775.900 458.570 1890.640 ;
        RECT 462.470 1775.900 548.570 1890.640 ;
        RECT 552.470 1775.900 638.570 1890.640 ;
        RECT 642.470 1775.900 728.570 1890.640 ;
        RECT 732.470 1775.900 818.570 1890.640 ;
        RECT 12.470 1774.080 818.570 1775.900 ;
        RECT 15.970 1343.040 818.570 1774.080 ;
        RECT 12.470 1340.640 818.570 1343.040 ;
        RECT 12.470 1225.900 98.570 1340.640 ;
        RECT 102.470 1225.900 188.570 1340.640 ;
        RECT 192.470 1225.900 278.570 1340.640 ;
        RECT 282.470 1225.900 368.570 1340.640 ;
        RECT 372.470 1225.900 458.570 1340.640 ;
        RECT 462.470 1225.900 548.570 1340.640 ;
        RECT 552.470 1225.900 638.570 1340.640 ;
        RECT 642.470 1225.900 728.570 1340.640 ;
        RECT 732.470 1225.900 818.570 1340.640 ;
        RECT 12.470 1224.640 818.570 1225.900 ;
        RECT 15.970 793.600 818.570 1224.640 ;
        RECT 12.470 790.640 818.570 793.600 ;
        RECT 12.470 675.900 98.570 790.640 ;
        RECT 102.470 675.900 188.570 790.640 ;
        RECT 192.470 675.900 278.570 790.640 ;
        RECT 282.470 675.900 368.570 790.640 ;
        RECT 372.470 675.900 458.570 790.640 ;
        RECT 462.470 675.900 548.570 790.640 ;
        RECT 552.470 675.900 638.570 790.640 ;
        RECT 642.470 675.900 728.570 790.640 ;
        RECT 732.470 675.900 818.570 790.640 ;
        RECT 12.470 675.200 818.570 675.900 ;
        RECT 15.970 244.160 818.570 675.200 ;
        RECT 12.470 240.640 818.570 244.160 ;
        RECT 12.470 10.240 98.570 240.640 ;
        RECT 102.470 10.240 188.570 240.640 ;
        RECT 192.470 10.240 278.570 240.640 ;
        RECT 282.470 10.240 368.570 240.640 ;
        RECT 372.470 10.240 458.570 240.640 ;
        RECT 462.470 10.240 548.570 240.640 ;
        RECT 552.470 10.240 638.570 240.640 ;
        RECT 642.470 10.240 728.570 240.640 ;
        RECT 732.470 10.240 818.570 240.640 ;
        RECT 822.470 10.240 908.570 2939.680 ;
        RECT 912.470 10.240 998.570 2940.640 ;
        RECT 1002.470 10.240 1088.570 2940.640 ;
        RECT 1092.470 10.240 1178.570 2940.640 ;
        RECT 1182.470 10.240 1268.570 2940.640 ;
        RECT 1272.470 10.240 1358.570 2940.640 ;
        RECT 1362.470 10.240 1448.570 2940.640 ;
        RECT 1452.470 10.240 1538.570 2940.640 ;
        RECT 1542.470 10.240 1628.570 2940.640 ;
        RECT 1632.470 2940.640 2258.570 2942.400 ;
        RECT 1632.470 10.240 1718.570 2940.640 ;
        RECT 1722.470 10.240 1808.570 2940.640 ;
        RECT 1812.470 10.240 1898.570 2940.640 ;
        RECT 1902.470 10.240 1988.570 2940.640 ;
        RECT 1992.470 2325.900 2078.570 2940.640 ;
        RECT 2082.470 2325.900 2168.570 2940.640 ;
        RECT 2172.470 2325.900 2258.570 2940.640 ;
        RECT 2262.470 2325.900 2348.570 3467.145 ;
        RECT 2352.470 2325.900 2438.570 3467.145 ;
        RECT 2442.470 2325.900 2528.570 3467.145 ;
        RECT 2532.470 2325.900 2618.570 3467.145 ;
        RECT 2622.470 2325.900 2708.570 3467.145 ;
        RECT 2712.470 2325.900 2798.570 3467.145 ;
        RECT 2802.470 2326.240 2870.105 3467.145 ;
        RECT 1992.470 1890.640 2798.570 2325.900 ;
        RECT 1992.470 1775.900 2078.570 1890.640 ;
        RECT 2082.470 1775.900 2168.570 1890.640 ;
        RECT 2172.470 1775.900 2258.570 1890.640 ;
        RECT 2262.470 1775.900 2348.570 1890.640 ;
        RECT 2352.470 1775.900 2438.570 1890.640 ;
        RECT 2442.470 1775.900 2528.570 1890.640 ;
        RECT 2532.470 1775.900 2618.570 1890.640 ;
        RECT 2622.470 1775.900 2708.570 1890.640 ;
        RECT 2712.470 1775.900 2798.570 1890.640 ;
        RECT 2805.970 1889.760 2870.105 2326.240 ;
        RECT 2802.470 1776.800 2870.105 1889.760 ;
        RECT 1992.470 1340.640 2798.570 1775.900 ;
        RECT 1992.470 1225.900 2078.570 1340.640 ;
        RECT 2082.470 1225.900 2168.570 1340.640 ;
        RECT 2172.470 1225.900 2258.570 1340.640 ;
        RECT 2262.470 1225.900 2348.570 1340.640 ;
        RECT 2352.470 1225.900 2438.570 1340.640 ;
        RECT 2442.470 1225.900 2528.570 1340.640 ;
        RECT 2532.470 1225.900 2618.570 1340.640 ;
        RECT 2622.470 1225.900 2708.570 1340.640 ;
        RECT 2712.470 1225.900 2798.570 1340.640 ;
        RECT 2805.970 1340.320 2870.105 1776.800 ;
        RECT 1992.470 790.640 2798.570 1225.900 ;
        RECT 2802.470 1221.920 2870.105 1340.320 ;
        RECT 2805.970 790.880 2870.105 1221.920 ;
        RECT 1992.470 675.900 2078.570 790.640 ;
        RECT 2082.470 675.900 2168.570 790.640 ;
        RECT 2172.470 675.900 2258.570 790.640 ;
        RECT 2262.470 675.900 2348.570 790.640 ;
        RECT 2352.470 675.900 2438.570 790.640 ;
        RECT 2442.470 675.900 2528.570 790.640 ;
        RECT 2532.470 675.900 2618.570 790.640 ;
        RECT 2622.470 675.900 2708.570 790.640 ;
        RECT 2712.470 675.900 2798.570 790.640 ;
        RECT 1992.470 240.640 2798.570 675.900 ;
        RECT 2802.470 672.480 2870.105 790.880 ;
        RECT 2805.970 241.440 2870.105 672.480 ;
        RECT 1992.470 10.240 2078.570 240.640 ;
        RECT 2082.470 10.240 2168.570 240.640 ;
        RECT 2172.470 10.240 2258.570 240.640 ;
        RECT 2262.470 10.240 2348.570 240.640 ;
        RECT 2352.470 10.240 2438.570 240.640 ;
        RECT 2442.470 10.240 2528.570 240.640 ;
        RECT 2532.470 10.240 2618.570 240.640 ;
        RECT 2622.470 10.240 2708.570 240.640 ;
        RECT 2712.470 10.240 2798.570 240.640 ;
        RECT 2802.470 10.240 2870.105 241.440 ;
        RECT 7.230 2.895 2870.105 10.240 ;
      LAYER met5 ;
        RECT 7.020 2988.790 2844.060 2997.900 ;
        RECT 7.020 2898.790 2844.060 2982.490 ;
        RECT 7.020 2808.790 2844.060 2892.490 ;
        RECT 7.020 2718.790 2844.060 2802.490 ;
        RECT 7.020 2628.790 2844.060 2712.490 ;
        RECT 7.020 2538.790 2844.060 2622.490 ;
        RECT 7.020 2448.790 2844.060 2532.490 ;
        RECT 7.020 2358.790 2844.060 2442.490 ;
        RECT 7.020 2268.790 2844.060 2352.490 ;
        RECT 7.020 2178.790 2844.060 2262.490 ;
        RECT 7.020 2088.790 2844.060 2172.490 ;
        RECT 7.020 1998.790 2844.060 2082.490 ;
        RECT 7.020 1908.790 2844.060 1992.490 ;
        RECT 7.020 1823.490 2844.060 1902.490 ;
        RECT 7.020 1818.790 97.370 1823.490 ;
        RECT 643.670 1818.790 2077.370 1823.490 ;
        RECT 2623.670 1818.790 2844.060 1823.490 ;
        RECT 7.020 1728.790 2844.060 1812.490 ;
        RECT 7.020 1638.790 2844.060 1722.490 ;
        RECT 7.020 1548.790 2844.060 1632.490 ;
        RECT 7.020 1458.790 2844.060 1542.490 ;
        RECT 7.020 1368.790 2844.060 1452.490 ;
        RECT 7.020 1283.490 2844.060 1362.490 ;
        RECT 7.020 1278.790 97.370 1283.490 ;
        RECT 643.670 1278.790 2077.370 1283.490 ;
        RECT 2623.670 1278.790 2844.060 1283.490 ;
        RECT 7.020 1188.790 2844.060 1272.490 ;
        RECT 7.020 1098.790 2844.060 1182.490 ;
        RECT 7.020 1008.790 2844.060 1092.490 ;
        RECT 7.020 918.790 2844.060 1002.490 ;
        RECT 7.020 828.790 2844.060 912.490 ;
        RECT 7.020 738.790 2844.060 822.490 ;
        RECT 7.020 727.790 97.370 732.490 ;
        RECT 643.670 727.790 2077.370 732.490 ;
        RECT 2623.670 727.790 2844.060 732.490 ;
        RECT 7.020 648.790 2844.060 727.790 ;
        RECT 7.020 558.790 2844.060 642.490 ;
        RECT 7.020 468.790 2844.060 552.490 ;
        RECT 7.020 378.790 2844.060 462.490 ;
        RECT 7.020 288.790 2844.060 372.490 ;
        RECT 7.020 198.790 2844.060 282.490 ;
        RECT 7.020 108.790 2844.060 192.490 ;
        RECT 7.020 18.790 2844.060 102.490 ;
        RECT 7.020 7.700 2844.060 12.490 ;
  END
END user_project_wrapper1
END LIBRARY

